netcdf weather {
dimensions:
    time = 3 ;
variables:
    float time(time) ;
        time:units = "days since 2014-01-01 00:00" ;
    float temp(time) ;
        temp:units = "degrees_c" ;
    float rainfall(time) ;
        rainfall:units = "mm" ;
// global attributes:
    :comment = "Created as an exercise" ;
data:
 time = 0, 0.5, 1 ;
 temp = 2.34, 6.7, -1.34 ;
 rainfall = 4.45, 8.34, 10.25 ;
}